interface chromite_intf(input bit CLK,RST_N);
endinterface

